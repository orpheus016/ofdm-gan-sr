//==============================================================================
// Tanh Activation Module
//
// Implements tanh(x) using piecewise linear approximation (PLAN)
//
// tanh(x) ≈ 
//   x                     if |x| < 1
//   sign(x) * (1 - 1/|x|) if 1 <= |x| < 4
//   sign(x)               if |x| >= 4
//
// Or using LUT for better accuracy
//
// Fixed-Point: Q8.8 (16-bit signed)
//==============================================================================

module activation_tanh #(
    parameter DATA_WIDTH = 16,             // Q8.8 format
    parameter USE_LUT    = 1,              // 0: PLAN approx, 1: LUT
    parameter LUT_DEPTH  = 256,            // LUT entries (8-bit address)
    parameter PIPELINED  = 1
)(
    input  wire                         clk,
    input  wire                         rst_n,
    input  wire signed [DATA_WIDTH-1:0] data_in,
    input  wire                         valid_in,
    output wire signed [DATA_WIDTH-1:0] data_out,
    output wire                         valid_out
);

    //--------------------------------------------------------------------------
    // LUT-based Tanh
    //--------------------------------------------------------------------------
    generate
        if (USE_LUT) begin : gen_lut
            
            // LUT stores tanh values for positive inputs [0, 4) in Q8.8
            // Address: input[11:4] gives 256 entries for range [0, 4)
            // Negative inputs: tanh(-x) = -tanh(x)
            
            reg [DATA_WIDTH-1:0] tanh_lut [0:LUT_DEPTH-1];
            
            // Initialize LUT (tanh values)
            // tanh(x) where x = addr * 4/256 = addr/64
            initial begin
                // Generated using: round(tanh(i/64) * 256) for Q8.8
                tanh_lut[0]   = 16'h0000;  // tanh(0.000) = 0.000
                tanh_lut[1]   = 16'h0004;  // tanh(0.016) = 0.016
                tanh_lut[2]   = 16'h0008;  // tanh(0.031) = 0.031
                tanh_lut[3]   = 16'h000C;  // tanh(0.047) = 0.047
                tanh_lut[4]   = 16'h0010;  // tanh(0.063) = 0.063
                tanh_lut[5]   = 16'h0014;  // tanh(0.078) = 0.078
                tanh_lut[6]   = 16'h0018;  // tanh(0.094) = 0.094
                tanh_lut[7]   = 16'h001C;  // tanh(0.109) = 0.109
                tanh_lut[8]   = 16'h0020;  // tanh(0.125) = 0.124
                tanh_lut[9]   = 16'h0024;  // tanh(0.141) = 0.140
                tanh_lut[10]  = 16'h0028;  // tanh(0.156) = 0.155
                tanh_lut[11]  = 16'h002C;  // tanh(0.172) = 0.170
                tanh_lut[12]  = 16'h002F;  // tanh(0.188) = 0.186
                tanh_lut[13]  = 16'h0033;  // tanh(0.203) = 0.200
                tanh_lut[14]  = 16'h0037;  // tanh(0.219) = 0.215
                tanh_lut[15]  = 16'h003A;  // tanh(0.234) = 0.229
                tanh_lut[16]  = 16'h003E;  // tanh(0.250) = 0.244
                tanh_lut[17]  = 16'h0041;  // tanh(0.266) = 0.258
                tanh_lut[18]  = 16'h0045;  // tanh(0.281) = 0.272
                tanh_lut[19]  = 16'h0048;  // tanh(0.297) = 0.286
                tanh_lut[20]  = 16'h004B;  // tanh(0.313) = 0.300
                tanh_lut[21]  = 16'h004E;  // tanh(0.328) = 0.313
                tanh_lut[22]  = 16'h0052;  // tanh(0.344) = 0.326
                tanh_lut[23]  = 16'h0055;  // tanh(0.359) = 0.339
                tanh_lut[24]  = 16'h0058;  // tanh(0.375) = 0.352
                tanh_lut[25]  = 16'h005B;  // tanh(0.391) = 0.365
                tanh_lut[26]  = 16'h005D;  // tanh(0.406) = 0.377
                tanh_lut[27]  = 16'h0060;  // tanh(0.422) = 0.389
                tanh_lut[28]  = 16'h0063;  // tanh(0.438) = 0.401
                tanh_lut[29]  = 16'h0065;  // tanh(0.453) = 0.412
                tanh_lut[30]  = 16'h0068;  // tanh(0.469) = 0.424
                tanh_lut[31]  = 16'h006A;  // tanh(0.484) = 0.435
                // ... Continue pattern for saturation region
                // Simplified: fill remaining with interpolation to 1.0
                tanh_lut[32]  = 16'h006D;
                tanh_lut[48]  = 16'h0080;
                tanh_lut[64]  = 16'h0092;  // tanh(1.0) ≈ 0.762
                tanh_lut[80]  = 16'h00A1;
                tanh_lut[96]  = 16'h00AC;  // tanh(1.5) ≈ 0.905
                tanh_lut[112] = 16'h00B4;
                tanh_lut[128] = 16'h00BA;  // tanh(2.0) ≈ 0.964
                tanh_lut[144] = 16'h00BE;
                tanh_lut[160] = 16'h00C1;
                tanh_lut[176] = 16'h00C4;
                tanh_lut[192] = 16'h00C6;  // tanh(3.0) ≈ 0.995
                tanh_lut[208] = 16'h00C8;
                tanh_lut[224] = 16'h00C9;
                tanh_lut[240] = 16'h00CA;
                tanh_lut[255] = 16'h00CB;  // tanh(4.0) ≈ 0.999
                
                // Fill intermediate values (linear interpolation in synthesis)
                // In real implementation, generate full table
            end
            
            // Logic
            wire is_negative;
            wire [DATA_WIDTH-1:0] abs_input;
            wire [7:0] lut_addr;
            wire saturated;
            reg [DATA_WIDTH-1:0] lut_value;
            wire signed [DATA_WIDTH-1:0] result;
            
            assign is_negative = data_in[DATA_WIDTH-1];
            assign abs_input = is_negative ? (~data_in + 1) : data_in;
            
            // Address: abs_input / 16 (shift right by 4), saturate to 255
            assign saturated = (abs_input[DATA_WIDTH-1:12] != 0);  // |x| >= 16
            assign lut_addr = saturated ? 8'hFF : abs_input[11:4];
            
            // LUT lookup
            always @(*) begin
                lut_value = tanh_lut[lut_addr];
            end
            
            // Apply sign
            assign result = is_negative ? (~lut_value + 1) : lut_value;
            
            // Pipeline register
            if (PIPELINED) begin : gen_pipe
                reg signed [DATA_WIDTH-1:0] data_out_reg;
                reg valid_out_reg;
                
                always @(posedge clk or negedge rst_n) begin
                    if (!rst_n) begin
                        data_out_reg <= 0;
                        valid_out_reg <= 1'b0;
                    end else begin
                        data_out_reg <= result;
                        valid_out_reg <= valid_in;
                    end
                end
                
                assign data_out = data_out_reg;
                assign valid_out = valid_out_reg;
            end else begin : gen_comb
                assign data_out = result;
                assign valid_out = valid_in;
            end
            
        end else begin : gen_plan
            //------------------------------------------------------------------
            // Piecewise Linear Approximation (PLAN)
            //------------------------------------------------------------------
            wire is_negative;
            wire [DATA_WIDTH-1:0] abs_input;
            wire signed [DATA_WIDTH-1:0] result;
            
            assign is_negative = data_in[DATA_WIDTH-1];
            assign abs_input = is_negative ? (~data_in + 1) : data_in;
            
            // Thresholds in Q8.8
            localparam [DATA_WIDTH-1:0] THRESH_1 = 16'h0100;  // 1.0
            localparam [DATA_WIDTH-1:0] THRESH_4 = 16'h0400;  // 4.0
            localparam [DATA_WIDTH-1:0] ONE      = 16'h0100;  // 1.0
            
            wire [DATA_WIDTH-1:0] plan_result;
            
            // PLAN segments
            assign plan_result = 
                (abs_input < THRESH_1) ? abs_input :                    // Linear region
                (abs_input < THRESH_4) ? (ONE - (ONE / abs_input)) :    // Saturation region (approx)
                ONE;                                                     // Saturated
            
            assign result = is_negative ? (~plan_result + 1) : plan_result;
            
            if (PIPELINED) begin : gen_pipe_plan
                reg signed [DATA_WIDTH-1:0] data_out_reg;
                reg valid_out_reg;
                
                always @(posedge clk or negedge rst_n) begin
                    if (!rst_n) begin
                        data_out_reg <= 0;
                        valid_out_reg <= 1'b0;
                    end else begin
                        data_out_reg <= result;
                        valid_out_reg <= valid_in;
                    end
                end
                
                assign data_out = data_out_reg;
                assign valid_out = valid_out_reg;
            end else begin : gen_comb_plan
                assign data_out = result;
                assign valid_out = valid_in;
            end
        end
    endgenerate

endmodule
